module decrypt1_stimulus;
wire [1:64]cip_text2;
reg [1:64]cip_text1;
reg [1:48]key1,key2,key3,key4,key5,key6,key7,key8,key9,key10,key11,key12,key13,key14,key15,key16;
decrypt decryption1(cip_text2,cip_text1,key1,key2,key3,key4,key5,key6,key7,key8,key9,key10,key11,key12,key13,key14,key15,key16);
initial
begin
$monitor("cip_text2=%b,cip_text1=%b",cip_text2,cip_text1);
cip_text1=64'b10000101_11101000_00010011_01010100_00001111_00001010_10110100_00000101;
key1=48'b000110_110000_001011_101111_111111_000111_000001_110010;
key2=48'b011110_011010_111011_011001_110110_111100_100111_100101;
key3=48'b010101_011111_110010_001010_010000_101100_111110_011001;
key4=48'b011100_101010_110111_010110_110110_110011_010100_011101;
key5=48'b011111_001110_110000_000111_111010_110101_001110_101000;
key6=48'b011000_111010_010100_111110_010100_000111_101100_101111;
key7=48'b111011_001000_010010_110111_111101_100001_100010_111100;
key8=48'b111101_111000_101000_111010_110000_010011_101111_111011;
key9=48'b111000_001101_101111_101011_111011_011110_011110_000001;
key10=48'b101100_011111_001101_000111_101110_100100_011001_001111;
key11=48'b001000_010101_111111_010011_110111_101101_001110_000110;
key12=48'b011101_010111_000111_110101_100101_000110_011111_101001;
key13=48'b100101_111100_010111_010001_111110_101011_101001_000001;
key14=48'b010111_110100_001110_110111_111100_101110_011100_111010;
key15=48'b101111_111001_000110_001101_001111_010011_111100_001010;
key16=48'b110010_110011_110110_001011_000011_100001_011111_110101;
end

endmodule
